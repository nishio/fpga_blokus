module main();
endmodule